module psl_tb;

endmodule : psl_tb




module dut_top (
);



endmodule
